`timescale 1ns/100ps/*Time Unit(ns)/Precision*/

`define width 8
`define cwidth 4

`define no_of_trans 8;
