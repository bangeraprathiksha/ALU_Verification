
`define width 8
`define cwidth 4

`define no_of_trans 2000
